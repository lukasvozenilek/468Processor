module Decoder4_16 (out, in);
	input [3:0] in;
	output reg [15:0] out;

	always@ (*)
	begin
		case(in)
			4'd0: out = 16'b0000000000000001;
			4'd1: out = 16'b0000000000000010;
			4'd2: out = 16'b0000000000000100;
			4'd3: out = 16'b0000000000001000;
			4'd4: out = 16'b0000000000010000;
			4'd5: out = 16'b0000000000100000;
			4'd6: out = 16'b0000000001000000;
			4'd7: out = 16'b0000000010000000;
			4'd8: out = 16'b0000000100000000;
			4'd9: out = 16'b0000001000000000;
			4'd10:out = 16'b0000010000000000;
			4'd11:out = 16'b0000100000000000;
			4'd12:out = 16'b0001000000000000;
			4'd13:out = 16'b0010000000000000;
			4'd14:out = 16'b0100000000000000;
			4'd15:out = 16'b1000000000000000;
			default: out = 0;
		endcase
	end
endmodule  